module test();

    initial begin 
        $display("hello");
    end
endmodule
